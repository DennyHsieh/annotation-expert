BZh91AY&SY�l� �߹Xy����߰���� 
 � ``	~K�J��t%$IJ��2dшi����4ɈMi�0� ��F�   �  2dшi����4ɈMi�0��A4�4� L&  #hɈ4�$�4L��4)����� z����� � ��jb$�ҏQ���~� dh m@57��C�U
E@�����(�(�$(���(į�J�H\�E�U4�L��$�IRN��s�Q0H#����L�:����_��;��go����ݻ��{�B��n��W�R���ג������\z>��"����:A�%?���7)��j3L�k��������P�
"�,υq�3�{"�ڛ&����/j+��ִ��6�-6�icE�Y�rP���'U-Un�/�5�ѯQ����pO ܒ�q��5&��m�Bŋ36�al�@�3\1Oc�@�A/�6����)�]&�'T�0�үK�-oD�q������̫�����5����v���C�;���D@QP�?.]>N��r=�"fT��8p�Pbվ��q8�77����A�r=�9^�Ȱͨ��f$��3$T2�K�F>�X��@ԃ�Mh'$�nP���`,0唁�$c	֕�҃j]T*����c�#X�sX��Ďe􈲶��C��P:u�Xuɧm��}LmX�Ր��V*�-`�%y�[����;P�K4�
A�Gsu���W�� ��i}A��O�؈lmV߆��z�a:Ҿ<�(�D=U�59VZ]?HN�l����|nJ����d޲����_u)����me����š̦0���C�!F�HSjm؅�S�kM�(���d�H�V�����[xT(�4�ڊ7l�Y=B���!Q�tU�#X�L���E��͍��t/	 ��)�x7]�5��D���!!5Ip��Y0*(mE�u�)�%q�7��O~�#��[M��[>����$2L%$�I$�I1$��D�����+�JD�u�咒�qIIIHN�D��p��4�	
����
�ZB����%�D̒�P�J�RZ�a�*�([Z�`eD���!(��A��A%����RRhH�&	@��K1w�BH�B$ (H��|!ZS���M1��c�̻�rrVD�`���
���9�"d�SV�}	ݒc�(�0NT��YL�J&d��5�'�]i�d�����'�'�:r$�T=�Ѝ�M#�"[�MY&B��֬JD��o�`�`	��zL�� ��I&e�WaE��� �)�.�~�IIOJ`�PR�5����	�8���B�N.�ҕJ@�<ə;�?�.����b�	�qZR.��� �j���.1G�:�5��`�1b�(��ҝ&A����%�h��#��e:MF sM���%ՠ8	�T�v�zO.	�¤*�&ѥ<��ԗ)Λӊ`���::D���K� j�pHM�^	�	���橐x	a7�kK�����8UC��:dt/�lSA/K�j��#�W�j�v�I�����HC�)
mK)��u�k��H�J"u�kl�N``K&�&BPU`V�x��h }唑�XƣA�������ح�H&� �h��KY"�	��e���=�ؔ(M�&J��%zSP�,�>)��p�O�M�Y�z�p�7�N�y�z<��=���M	p"hJMȏ:�b��ޝ
��],'�И	�`�:���i@�Ad	� t�74V�u�$��X�r���֮t���!<��od�D�%F�2��Y1�P%���PrN��H4���9�Rɀ%'2`�.� �)TCN�b'�$���I#dؖ��K#��Or%)m��$W�����聓؂����<��H�
��� 