BZh91AY&SYWa/8 ߹xy����߰���� 
 � ``	�yg�:�@ =��4R�(IJQO�1�L�ɠ  4�  �&�M��@�    �F�142a4��4ɡ�@a&�� � 4h       "�4A�hR==<�����(�=A��z�=AQ56�i=O � @ � [�R#�%* l
�z�_��Ѫ�2@&� $�0N�����X��B%#	��
��YRk@V����x"41P�"$�K��sW!�c�P�u��(R]��g���f�_&��M%�� �B�nBD�H'�IM��c�Č"W�Q�ŌN��_+�4�e�C�a@�=��n��hi�ӎ[��}'�KQEQ*�vS���ק7��iqն�wt���S8��5+�Ks��'�~J/hVEQ;�� �7��t��+^� q.a�[F�&X����W��8(���s�՘Y�fjJD�S�0���u-�QP��&L�F+h��(^\\`^��U��Vb\�����=_�:��L;��'"@`'ߋ�ǻ�^� ��+�Wd��VwƗ>��q^�`.��m����D�;��
�ɣ�8[~jT�c�^rI�Wx$�ZGza�uj�3G�����N��	�(�Ȑ�h������jU6��ʌ��m�Q�eTҎK@�Tm�3�+F���I����v<��UWQ�&/�%Z��@=�-Kl`��q**E16s!����]HuA|��9�O�5V��u2�n�	սH�SYq}F�.�w��|�,p��]�U�o2b7ԵZ�Q�Q6�N�.��2�S+�"�6��֫9	�J�4sG��
�9�h�b��t٥���D�[hK�̊rۆ�ƙ6��b�F_Ȳ��jŪ�L-:p6�l�}ڂw���<Z���f�Y��V�Jh�}�E�gf�`�틭[k��.n"ؽB+�W�J���%�%��ڸ��2�iY*'�>�8u8��� ��"�"�"$]ꢊ
�*��� �����C���VV�h��dddRt	��f�MZ��,��ʘJ�bf(�(=�h�eR�1��F	��Q����2�*P�beTU��A�D�(I�d��$
R`��646��!c �0��f*�,Y 
I��0�7nO</?�si��d�Fn&#j�m�~3�P;��$�8ӡu�-�Ÿ����4�zF����G��7н`\��_{���b��6�^hPN5H펑�G��\�ĉp��AT$ �y�̼�C�:�P!`��(H�A;�X���p���C�B�v������@��
M��V�)i HC�mP��@�����Di+`4���Kw��<�p��&����F���m��9��?2Im�wV(���IF@�dj0�0<�쓎�u|��.0r�!��F �@���o����\��;A�N�q*����.�28�`��Ph8>`�OQ�TsjF���eaƄ���>A�z�?�6{��a�7#YP�������h�8;���`;A�p�����`v��(���s#y>7.å�肫�D=(p9�߸|��4�u�Q�X�޷.�m4�DNA�GP�GM04��R�P�*���R�+�dc�f��Q̡e�����T1���(BZ�Өx�I�����`��7��f�H�/�=�c�pP�C���8���m��X�)�w�R�/G� ��1@5(E�Ǫ:DCH�e���6��E�����Z����[Pe�D�Զ��Xλ�H��n(A�}�D.P��^M�����6-2�D*<��p��Z�JD�2@p� �����_��rG.��U@{F�S?V�BZ2��/���j:ƹEp3��H�t�`��[w�-�0`��`��7�A�����|o�.�p� ��^p