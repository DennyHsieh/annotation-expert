BZh91AY&SY.J �_�xy����߰���� 
 � ``	_=e��t�� ��v�Q!*IQO=A����    ��	�*jh h      d��dɄ� d4��&� M���SG����@b4� 2�M �I��56���iLe�ѧ��OQ��4ɑ�I#H�F���=C��=A���h4��������U
Q ��=�w�T�D�J
�� q`��S�`{�(����QL�ຫR��L8��{ 41�43�9M5K[Q�k��d[�x��o���G��c8��QH�'s�&z����S�a�L�3A��@�"���ӱ|�`�޸ZT;q��]um�P{!�1C�ǎkө��<�������g*aN=)8�����rT�rt�/x���z)+�E�gg��	�C*�M��Ri���0tg+^����
*,*%f��Me#m������:��W��	�f`�f
8�iD��$�L�q�ߏ��pp�����!HT�=���.߽�o�W���3pfM��`Ȩ�e4
�c�dC͏>o\�]&V�%���'py�l^�ֈ�Ӈ��3<$0z�����#`���m�ҖRRd#�L��	z���bd��bp���/0�JA�]T�Aǒ�CT�$괄Ƹ܂��h�s8�nDn�h�b��pf���܁��Z�ֵʜb�VZ��5�47]jC�R����5���Z�.8av$U�ddo�U���ںG%;��i�v�:j�WX�y��:x�j�a���xd��q ݄����^-Zf�v�V�PȢ�@;�4<�ȠcQ���,V\��.,bFw��Ubh4��O�E���+kYV�q����Z�{��xw���WO}*�˛����v0%ډ&��V����whejڲ|з/<:�C��� �@�0$11�窪���U��EI}Xu�>��\���İՁ�JH=C��*DU �C���v	�RD$Ht�^�*E$D"�^�(��IjJ!kR��l�D�H���$(R��f��(	Pd-5LEhTAd�*.	��<�-��Qe^���.�
lH��!&<��`� x�`�R�.nLtᆵѣ�ױ(e�\8L�`]}�����)�.��	@��'�C!����d��F��I"�oP�Z�NA�0l{`���әBIB$�=C�t��.�s ��B��7���q��P��X�vؓ!�I&)R�ѾI$�JǜA����7��S��٪KZ��q��.R`���b�$�A��		0��b<�0U-Py�
JH��0ha9����Rޯ�~E�LF�C�(�Y�^��\RD�3��:t$���4u�#�I� i���#�|�)v�`�)7��;�P���Ӡr����JÐ֍2!�˛4���_�S1!S4m���r� ��Ծ H�_�xA��VcUq��!��W �C�s��Ǿ0?(��qS9��GH���Ch6����1M��qM�E,  6FѤC�0R��Xh`�J�%b�b�\`>�1h�t����R�D�LSp�Gj��5��r�@��0���/�>�I��
2�M汸�@;�(���~�ĵKh�ޒB nP���Ԟ � {�fK��epK���CA�\�A�#�R�F푰�/A��ڡ	�=��P�BƻD�h�%u%eP�Ƌn�R��H8��q�5)%)u�X�� �&��\jL� SIfѺ6��<����[��#z�'�iMCMf#B�d9���<!p0�ϫ9� !�0�Z8�����5����)��rP�