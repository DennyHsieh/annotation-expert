BZh91AY&SYZ�A  ߹xy����߰���� 
 � ``	��ϼ�޲ ��Tl� �	
j����I�@b   b@  % M"�� @      ��2bh2d�i�2@i�C &��MD�OP  ��4�ѐ �@ MTJz)��&�C�0���  �� "���e4�5?T�z�����F���G�z�����t�,ȫh+}O%��q����V���2�K�	�a7H�C X�rB%��*�@c8ǒo(o���0�3�`B�-�B����)t�
ڎ���4�B���y�K�8
���MSc8DOPS �Or1F܀{�����Ѐ��F2�ۄwz�&��!��7,���4�,G��%�(#�H&vu�u��EǾ�4#�(��]�z)��)�MSK�����h[�ǵʘyƧ���o,h4��-9^ZpM�s�4(����@RW~�j�VS��� ⺇Z�dr�A�`iy8:trQ'#��1�bޟ0�'*D� -�$�åkk�o[�c]����nKm���+.{b	by����u��;D���9D�`�=_����T�]8
�P�Uк��
�[�Y,-+x�F�	XV���C���B�xtp�o­J�Lc��I6���kZR"�i����T@��	����R��!h������\ �mJ���ۊ��ʩ��D�t�ۆf�V��%��I����v<���U�i�/�%Z��@=�-KM�����0��I�J�����8��]�z�ɮ�z�;"yEI��GK��{vHN�Ԍ�6	Hh�?D�M����F+��c��b��"ddo���ʌ����u�vg����_�鴕ƵX?!<�]4f�h�к�Z2MLB9]��C[4�[��.З�K�����2ms&Ŋ��7�ee�.�X�[ȅ��p>Uh�|%�	�ۅ��<Z���f�q��V��� J;����������Й�l������[%�	͈*��Q*��h���t"��.�̭ZVO�>姂Q�y� ��P�"$D��UUH�*���,�7�����fo\ɭ�Ή�J%��T�K��<��U�U��n�.�%P�
	��b�-Ub$Q�b�(d*�(�tK���*��nA�D�(I��A(HG�#Q�eF� t��1D�H� �@�������})<�f����ݧP&я*�#ה���}�m��X2���;�*�J�X��ٴh���S%�vxG����m�/]��@07R_�\ӵ8�y;�:~��"m�3Đڡ �Ҏ+�`hx��:�
���+3E3K�r�1��'j������lk���� P�ԡ3�zT� dsT<��dd}Cp���-A�,�o���8�Rh�h�v��5A0H���vɽ&p?qDR0��"
꘡��'BVVL��35�31<3��ի�w�p��byp�1SA#��4<>�� �;��N�y*���r�]�(��-��s9(�6���1%fv��;Y���;��6�t�4���
ja�6��+�T\����;��240~ j�a�p�wf��e��:"� ~é�j6ݎʹJ6 �%x�߼5V"���Nbwf�NY�o�Ω8��6LErSBuI���rF)���pSD��V#I��2+&��hd��L�{�:��8��d�;���n)�fF��lAI���x��qR7Vr��ަ�]��q����������9�����4�b���l��'n9fb�Γ�7[�֛ʗ�����XP�<�z�j�*�R��(tZxG�j�� �!mP�n	������ƅ�;�F�:��w>b��^݀9s���Ѹ��U��D,:�s��LJD�2@��H�ar�)�l��ͳj��+��lM5+5>)�����V'�2�*9�Mg$��1����|�ÄZm�g��`P�0,"�Cx�����w����rE8P�Z�A