BZh91AY&SY�`0� �_�Xy���߰���� 
 � ``yf�@h�   �D�i��F�� ���  4�E     4   i�4�ɄM a4i� 	5����@�4 !�4 4 T4�ɓM1��d  �"�! S�h�&j�S��G�MmSL2���&4YQ �%� b!���D$1 �/|�0`LH�	�
d�=�V�
�~0� M8$�t��Roc	���}��������e5�j٤<�L���`CP!����A�B���Sib���t-���F#T̶�@z�"`%XF�@�P�#v��0ϟF���U�`�(�.�c=�:�+���:��kj70���l,���ej.���Q>D0*	m�۰�MiT��R���9B�rƢ��f�c7�4O)�!2�*8�䕺�?::o�sLͭ�(x(`/���ߔ��6�b� �	B�Q�@��4�	�n­LqI.P�)��T�}�h��4Sd��$C�*���
����H#�U�[���1͘����j$�$�K��s�)�E[��p�["X.
���f`�
�K��P�T`2��P$�qmPcZ���P�X��N����n�nƀ��ڧM�"h�
�J�GL���MT�q/E� ��RD��[��FgIA��cl��� @�3�58J��dl60�4��$ld2
�ap.,8pj�J�XzW2����K��`0,�ɻz��Zͽ	��9%h[1�����CH!��q2����TE�a6�˛i�|�Ҵ��+��~1R�����)ޔU�,7LNׂh��E>Y�o,.qBn9A�p��p�7�d�/UQUV*��P�G��y2I�RF��HO5�PnE���+�ԫn��.誕PC���t	���RT��It�B�W4*S��	 ��hF��HIL���R�"��%��@T�TAdhH3��Cӆ}��zyv�p՛�
nH��xA��$>�]��MbKA��'J?�|6$��Z�$�'�좕H׭2J�@�Ԫj:�F)��}�?�w��y$*�T�<�gN���򛶊�O�IK�=����t�8�,}$}M���1A�V~���r�I�ؘ��鄔��L=H@4�h%/|2���ڝ�uDR�DpM|��HHHH�V��)�! aG� \R�� �JN��BJB}����G���U����,�㧟	K�d�&	���Mģ)ҙ�&� v�U�,%4p��wMbi %6��bm�5^��N�=��4��,0��1[֪�߂�|�S�Mp\�P�����9{���!8 ��$�$r���ȋV�ڌfM��Pw���|��R;R�r��&'c��08	k�����l�N�t��J���Ig�jH-��h�JBb�	`[�] |��At��.'�K$��r��@8p�n(��U�3 ��=)s��s��Ќ����&tޗN)	�&���rOZi:�*��
<���z��8 ��9���O�I��͒<�itr4�t�K H7d�j]�4R�ӊF��(�Bf7p颸J��d'N������V���=�Cڡ�CG�JD��5��5�	 ��1q9J`�
Y5�,��eh	o�] �}0�'�Ąq��y��e�^45�'�:8&P����؝� H@5fӒ~�~���� A�?��"�(H]0f�