BZh91AY&SY���% �_�Xy����߰���� 
 � ``	���O ) �C^�qI*@��h�de	�4=L424ё�4�F#M4	S�&�� @  �   p#	�!�@2 adɄ`!��IH�� 4       ��	꟪?J~�3OSS�2hh4@z �)��z�i�zA��  j�[R�
J��1 �6|bF�kF�	!5 L��>�`CE# Ȑ�%�X{�UV�Fb?1���(7E�B20(^ZV����0�$h*sJeG�֕E"�,�к@�V�B�)+|��9?}-��%�6�zT�v��,k��5,jiS�f~�t����$�	u�j�!U<� p��D�A�L�җmIo��
Eye�9^������2Ҝ�e�Sd�w�֠�LUfn.���T�O,4L��u�����&�Ryaf	����k՝'$s1�;��#�\$���饷j��� �[7�̲�EƖʴ�~]k�at�"%�r�+�Z������a:�[Vf���jD����M�9g�KZֵ��-kZ���y������(�*A^Ξ:��b�۹4�h#�]�[�[L�F9c��N5(� �ȹ��{/z�q�6��6�K�JN���ư�����	��[�Î[	��j��,BzH=���*L5\�CMZ����Q)���$g	
S;TK���[���;�b�G�$��u�I�6�Z�E����X%�튜�M3�e�F`a�ƭ��#40qJ�R�N�@M-+���G�l�����v�KM,1�k*��λ��:��>Ǎ��Z�|Ʈ�ֈ���6n�|a�����,,a��ef��[i��7X�mݦk��:�����i[m7
��&P�PI1�6`�b�%��x1�%E,a��An�aњw#,n�%�Lj�W$��y�Ι\3j[/��%q��k��ޫD���@6���D+��w�r3�}��Y��V�.�{d�d��Ғ(P�����Zvʃv��&a��hƻ9����lr�m
�p�������hWI�$F���m��}G|b"$]򪪢����H����:Ǵ!Ē#�ֲ5$Ѝ�##"âMF5�&�Ն�E�;7F�&VԸ��PA����kR��`4����H!*�̤ʔ�2�U�j�(E�N�K,��h29F����#F�l,�H�2*� ��,��]���^f���-�pY@!+��0
Dav}*�E45-K��<	�h�:q���~j����a�0� 0��hڙ/�1>ҝ�C�b!6J�����bW�-*X���':ͩ��09��Q=��)h�C�NV�,)(#f$��B$l������{j%j-[�7���ۮ"����Ǔ�\���E�|�YЈ��D*�,=��^�BQ��%,0�5�����K� 5�4��1B�@C,A)��I�tz����h7SЫ�J�<�V!w<2G���(. ��K�!��`�T`I���u���t��<"93�	R�r`�CU�N)���}�t�<�3�la�tr�Է0�D��D��Gj9d�\���k�Ҩ�ƅ�
�
SriMCD#�J�Ȩrظn0o�<�u�00�m0h*"-�V堡��FV�c�FR;l(X]��!!d��ƔHF��A� ȄRY�u8�QH���Q5@!�:��	�{G�t�Ru�C�u�H!��RPPl�X�G2��h�)�N��/�L��ARq 4B��a�≼_P}f#q<w�s�6���-�%�'NջAf��������: aw����!�QC �0zj��r�`�2΢�a�r�:R��LL��k�,�Rz�\^�7��HO6��\@{F��Ս��>Te�B[֡�*�fJ��p�G�pいNEX�#���`�h�p���q�n?�w$S�	
���P