BZh91AY&SYK�� _�xy���������� 
 � ``	��ϼ�Ѐ oC��kI%HTU����hi� hѠ  M2  P"(�M  �    ��2bh2d�i�2@i�C &��MD�OP4 hh�Ѡ h @h�I�F��j&�@z�4  ���"� MM�ʞ��=F��4����(XNz��J�A\
u��2�E�j��\�L� ���t�$1#��F0��UZ	^����1I�`:��L
ӄ�b/@@UY�!+��í;p���ݼi/<������.S�g�d�@܆��(2�f�E�#�%Ē ,�Lf)��7D ��5|j0/���@�>8�㓌EB�:�	�}N�-'��`L�EQ2�xS�[=wf�fwVԥ�B�K>��U0󦧕�ԯy�F�,�]�F	�6��
)�����Tc��3-�H�k�vZ���a$V�&Ru8(���X�Q�e"��ah�jw�� t]�J(�\�1�b�U
���Δ�S������?ׇ����v�cNQ��_r�" �oW�z  0Сjay8�j��Z�JD%`�b��t�~P�5)���#S)DƝ��$خ�$�f#�H�kY�U�"��y[ �A6�dHP�Hann#!SjP���kn*���SrZ
lT}�3�+F���I�e���y�-A*���1|�*�����Kw[�*�У�q*(E16s!����ފ�G�Y���'�T��Tt��G�d�鼑��ZyB˗�m���1�}l�Ћ��1x^�5��Z��Q�Q6�N��f{�$�W�EzlJ�2�9�O:2W7����
�9�0�1�5��$5�KE����	}���� ]�`�oTB�Sb�(��������jŪަ�U�l���2Jܣ�֖I���o���,�v���c��vf���gf�cK㋙m��ڹ��b�~�*��X�[��h%�9;Xx�VVO�>�xrt���O��"ȉ"�`���*������|�+�CU�24Y�Y��%�DI�L�%�i�g�
p����]�Swiv�v�����T�*�b�F	�����J@�]�.��]Ҩ
�nA�DI	�J�$B�BI�CFF��� \@�
�r*�,Y 
Gt Bw�t�'��c��L��Na��#���O��c�]��@ca�:SU�g��e�1��x���+a����E%�Wnm�gJt�)��u%�w�1�+�+*�(��13[���6ҴF�24�Wz_Y�l���7D�V�#�P�<'0<�l�@��
(L��J�@� �C�����8u��A��q������R�E�K�\���Q@4��&��@��U�H�N\��AiC��BJ2�#a���G�1s�G�t�4�k��l+T�(�$v)�훞�W<�`�<��N�ĕdg�;�^W�� �BE�>J��PB'Y��8��#VS��7�L�S:tO���+�&�ޕ4r�I�"��"�<:��`����5�0���\� ۘs��r�.� �l8�G",5*�V�rb$����E��=9�♰�ɡ8,�8�G-4�Do��":���6���,%b3�Fͦa_u�3�4̮�cFF>a�*Ge
\`dY0�iq��=�n�!���xdV���J�L�\ӊ�����ժ=��眇YEx�tL���a�n1<1ݘEϕ�:!۵��T��x
�r�`�i�M�Wv:nm��U=MD.	s�6P���-�e����K4f��Ƴt�2���X���;�2�2���@� ��r�`��+��-�:��Z�JD�2@f�:�"��s+qz(7p�}ra�3�L�~�:-{JbyS$�Q��9͇Q������}��\
�ţg�1���"�8�jvO��N�c����"�(H%�H� 