BZh91AY&SYd��� �_�Xy����߰���� 
 � ``�}���` 6���)RJB&SMjh��   4hM"P�=#j   ��h 2da�a4�h2hɐ�	5�jFF�dd 24h "��I�OdjOSOS@zA��4�2hh�� �)���A�m�hd �h4h i�
@��%D�b����A�E((�όN�
7�^p $�࿒�B+�!9dH%�<P�*����o�ߧN��xc��j�l��ڴh��V�K���
�K	��d(�u6�t����n��1��H�`���m��1d@̦`T*Z(�ey7nČ3�2��+.`�EIecʬ.��>��<���z�N��dYʕ�Q'щV0��LN/�xH>X>|�r�p�7�N:��L�&ѪJ{2��P���jRM��eʕ5��b�/ll?b��jBֈ��|1��r��<���F�uci���A�P�ͨ;?T�vM{fbbA�#��'�wW�Ү����T��w��*��`��¸� 	�d��_Pv;|���pMI%d;��H�b�HCZ�
�N���Fg�����a��m����L��p0f�{�����Ygf�m�X+��0������MU��Ì�HI'3 J!�����E�&�<�M��Y�G0r��\�/\�����.�]&MӦ�9,,Z�:k�9kF0pH��z�����JC�qu 4�us-"��x��k�5U�bI�
�h��hsC�au@�2FN����ȸ�|��
p�n Ќt6s����+�.vK�Dܠd�:���id�K��Rd�*w�a�#[G"u��NS�{Gaӿ3��{�+.m+qx��`4�I7N������[VO�#r��GK u�]A��u�)"0^r������F��N�z��2X���`|TIH�2�nJ2�t��U��J�*��yС%�$D& RH]�K��.��U"�ĩM�@H)X�(F��G$�)T�J��)E��4X�*�) 
I�A��Y��In�Jw��/ד�)bG�CϊDr�~a�%�;D��7si�u��G�Ȕg��{m�桄lП^>Z����� �(�P�G8��v�/W���O(&#�0����֦���E�Ehڑ�Lj!Y�s��t\
m��BLq鰴0S���ư#�^,z�I!V%6�(���%%>���Q�CU�R��+ۤN���k��&��;9��%q$���YM�]3L1
<F�`&�� JH˦l020���P�C������
���D����9�5	y-�߾��bJ�)�1^+�A������ �:�&uڌ� ��Œ��%@6�Ji���6��|�*�1�X!�Z����0v�(&�!i��knQ�N`�rMGqQ�DX���e܌(f<�$Dy@Cʽgb(q;����;��E^�#��]$Gh5�P�d�x7�]6�H�XЩ ���2��RFɪ�#�Ly�l�dv�K�/|��.�0���	`D��&����!��9@B;`�Gm1�a@?�|CPp�\�q%���i�`�%�A�k����=)�|���LR����(��`aA�M�!������[$���Tx����b֑P���$��`�I�b�5T��$.g.�W	��!4�֘]:�+�%��7��5�j9�2�$Į��l�$�r����0T�i#f�4���ȗD-�\ Byєt*��=t�|WeY��w����9@�54����.��T�a�Ó ����u��ֶ��]��BA����