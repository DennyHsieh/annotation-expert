BZh91AY&SYտVv (_�xy����߰���� 
 � ``	�yg�{z �:��l��Q1MS�I�7���@  @h  � �5H4� ##�   �A�F�142a4��4ɡ�@a&���� ��4# h i� "�B��50h���Ȁi�i��OP�D�z�i�Tڞ&�������z	���ʩ �(��	tó�$i�����.&0 I{�6�&���H��%��>8*�A������`�¯~��BЅHZ,��^s %.��[R5�{N"6�g]$��0����64D�
d�Os�f#M�;��v!pЈ��2�A��l�nP�)Q��z˩xʁd~M�SG�.�k�9-������$$�]	n��3�jb�ea���S���ƣ�ы-ɼp���x���с7M�Q���m��(�:p��^q�:֣#�p�+H�4Ĝ�ōaR�06���k�)�.��5�0��C/��\ �j�����+h�mC�#x���z8i4j��B�
 �������1WO �t ��A�ק�Y���quJP%a[ϵ�C�=K� �y�6F�6ɘ"D>2�<d�,� @���B����	���'���#B�R"�.X�E��"A�R��o4�����B�6Qt��}J��QsWU(��q�{a\nWn-�jP�aDR��mԡG� E �>��`����/��Stx�
D�d��F�Tt�wH��*��J�:��١X!��CX����L����i�X�XGf{�H��ZWww8pq��ھX�F�L��d*`HvBڬ+��"8:@�1�pt�XlX�����oX�'*�Mc��8�l����!q�m�:�!]�a�D���i�4���}i$y2�am�º����ڄ���X�qN�*�r��'��l�H�EƋ�a�t����,l9��ΘBz�R,��/!UUUAb��`A$��P�}�"��U��BU�k�D�$�&%���+)��m�B�*��K���!��
�)ULD̕
X&5	C!P��D���*B�EX��D�(I�� �E	@���h��l2�"����8+8�*�,X��!	��}	=�{M�i�B��<J�V�:��~�o�2���su��P����4g��r����9������v�����'ꡐ�h����#ң��D(��	 $^�q^������T]݊4A�OR���Q�`(~j�Q���pl J��J>�� �#�ܡ�큑���Ȉ����r�<�vDR�E3��#R[J	2̝�i(�L(�F�X�0��̈JJ���F�?����W��5�`}P�0�H�9MO�ܕ�7���N�q*���9X]�(��-���v�(�e�h��
;VQ��$j�����~�x����7�iP�ȦC�ɘ���$h]�Ps�9�H8o �
����c��v�r0Z����ܡ:W(  P�C�>P9���`z�����<]�9-��`�Gx�m�ìXê��4��ֲ�w�FVä����21���du(R�|`��|a�F����H�TY�?8�
��Gp(G849X:V`_�|a~!���s�"�N�ƀ�i�n��.��RX�����5NIPeXP�=��5��>0�뢇8%� �w(h2 �b�	F�9u����4.��258� `�\[,2�������ÉA�V��PP��k�G#�m1)L� f:M :A�����^i��D�cr4�����TSF�522��q/:�<#�&����9c(����������9�1�a�����i�v�����)�����