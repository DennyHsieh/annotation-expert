BZh91AY&SYԼ� _�xy����߰���� 
 � ``	���^*� �
�r�)PDQL��4ޤ�M  �@  (iD��4  4�  �F�142a4��4ɡ�@a&����24�4�Ʉ� � (�!�hJ7���ڣ�)�6�=@�A�P4�=A��i��2���g� @��@�����U-C"���E�j��\�LP I�0O-����$���A�����I@YI?!�
���^�F��Q(�`BMi��MB��}}vP���V�灋�|��4�9��D�
@;R܄C�ܐM����<�S�WF<�3�:�������3�`����S�,��A:s�s�H���IQEQ*�VS���7��iqն�wt���S8��5+�Ks��'x��UE�
�y�� �7��j�۷W$u��w���vi��s�RV�Ӓ�9�;8h�.�#D�eyq;�Dw�]�QPľ�Z���E�CB��S��&Y�%b%�pA,O���i�]L�	�˭�p ��0�o/���>%�@����-NK�.�͗V���{Q`��dC�0��~(P�E)���R����M���$��;��Y�D
�a �P�	�(�"B��C�7�ATڔ/*2�G��SJ9-�Q��3��X.��&oWw���Z�U]F�b��U��l���,M�����2��Sg2z_0����_,�Ns�*MU�:]L�۲Btޤe)�IB˧�oWk�F��d�p�݌U��L���Z�L�ʨ�{�]���h�JIl�Ȋ�ؕ��`�!<�]4f�h�к�[�$�t`�n܄rՎ�C[4�[��+p��$+K��Æ�ƙ6��b�F_Ȳ��jŪ�L-9�ڙ��Kj	�P�C�t�OWu�#{�g��V�Bh�;�B�7A!޺A�틙m��x�sq��_h*��X�[���-MF��ݸ�ej��}�3����;@�w��DH�9Q`��������V�|w�zFEm>�����%�DI�&"�x�1㲛YV�T.ҩ���Q�Px��*P�Ub$Q�L*�A�-���.��]Ҩ���H"��6J,h�$�G ё�lA��
0d2�D�Ȫ �d�)&b ���a��z;�Y�.�>^0&#uG��;��wCHI�q�Z�Z��1��UhP�v��Ə�o�z������D\0�s�d6('�CX���G���Gʉh��AT$ �x#�}����C��]�T$h� �������y_�P�� �r��� J�-E	��� H��6(ut@����҈�V�k��:����ݤ��*�q��(6� b=��8!�H�%�2A�kR�nD!%0��0�8H��'z��}a�W`;W1��F �@���+�3y���.@�x��OȢ�|�����Gj�k�����8�](��"8���q�#R<��0�>e�G~�5�:��k��E5��;�9�֍L� 6�1��v��P��D89r9����r'm����A̻ Uv�bN�7�a��b<r,�ظ��n0P�Q:��8�`8ꎰjD Z��+EC��[��+p���4�P����} b��q�#`>PkI��o6���R6T:�B8AC�7��f��6�[�mìpP�C��Ѡ8���l��.��R�޽�������a@7(B#�;DC@��@�)p�
(o����� 1�4G����ڋQ
��y!���P��=�\h��� vv���Q���k��`=7��#y�Z�%"I� �s8paeR�Z.�F��&��V� ?8Ԋf���A��#(ނ��c�k��5WC>#�h���r�.����7�A�n���|_�����H�
���`